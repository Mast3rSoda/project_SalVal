module flashing_diode_0_25s_board(
	input CLOCK_50,
	output [7:0] LEDR);
	
	flashing_diode_0_25s_board(CLOCK_50,LEDR);
	
endmodule