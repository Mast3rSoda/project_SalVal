module subtract_10_4_bits(
	input [3:0]x,
	output [3:0]A);
		
		assign A = x - 10;
	
endmodule