module circuitB(
	input [4:0]x,
	output [3:0]A);
		
		assign A = x - 10;
	
endmodule